module Project2(
input  [9:0] SW,
input  [3:0] KEY,
input  CLOCK_50,
input  FPGA_RESET_N,
output [9:0] LEDR,
output [6:0] HEX0,
output [6:0] HEX1,
output [6:0] HEX2,
output [6:0] HEX3
);
parameter DBITS                 = 32;
parameter INST_SIZE             = 32'd4;
parameter INST_BIT_WIDTH        = 32;
parameter START_PC              = 32'h40;
parameter REG_INDEX_BIT_WIDTH   = 4;
parameter ADDR_KEY              = 32'hF0000010;
parameter ADDR_SW               = 32'hF0000014;
parameter ADDR_HEX              = 32'hF0000000;
parameter ADDR_LEDR             = 32'hF0000004;
parameter ADDR_LEDG             = 32'hF0000008;

parameter IMEM_INIT_FILE        = "Sorter2.mif";
parameter IMEM_ADDR_BIT_WIDTH   = 11;
parameter IMEM_DATA_BIT_WIDTH   = INST_BIT_WIDTH;
parameter IMEM_PC_BITS_HI       = IMEM_ADDR_BIT_WIDTH + 2;
parameter IMEM_PC_BITS_LO       = 2;

parameter DMEMADDRBITS          = 13;
parameter DMEMWORDBITS          = 2;
parameter DMEMWORDS             = 2048;

// parameter OP1_ALUR              = 4'b0000;
// parameter OP1_ALUI              = 4'b1000;
// parameter OP1_CMPR              = 4'b0010;
// parameter OP1_CMPI              = 4'b1010;
// parameter OP1_BCOND             = 4'b0110;
// parameter OP1_SW                = 4'b0101;
// parameter OP1_LW                = 4'b1001;
// parameter OP1_JAL               = 4'b1011;

// Add parameters for various secondary opcode values

//PLL, clock generation, and reset generation
wire clk, lock;
//Pll pll(.inclk0(CLOCK_50), .c0(clk), .locked(lock));
PLL	PLL_inst (
    .refclk (CLOCK_50),
    .rst(!FPGA_RESET_N),
    .outclk_0 (clk),
    .locked (lock)
);

wire reset = ~lock;



// Put the code for getting opcode1, rd, rs, rt, imm, etc. here

// Create the registers

// Create ALU unit

// Put the code for data memory and I/O here

// KEYS, SWITCHES, HEXS, and LEDS are memory mapped IO

endmodule

